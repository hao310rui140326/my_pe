
module pow_m_0_75_fp16_encrypt_bb (

	input   clock,
	input   resetn,
	input   ivalid, 
	input   iready,
	output  ovalid, 
	output  oready,
	input   [15:0]  datain,
	output  [15:0]  dataout);
	

endmodule
