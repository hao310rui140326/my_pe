../pe_types.sv